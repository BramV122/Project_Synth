module Synth();


endmodule 